ENTITY entity_name IS
    PORT (
    port_1_name : mode data_type;
    ort_2_name : mode data_type;
    .......
    Port_n_name : mode data_type
    );
END entity_name;