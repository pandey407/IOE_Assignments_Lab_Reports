ENTITY entity_name IS  
    GENERIC (  
                  generic_1_name : data_type;  
                  generic_2_name : data_type;  
                   ........  
                  generic_n_name : data_type  
                   );  
 PORT (  
             port_1_name : mode data_type;  
              port_2_name : mode data_type;  
              ........  
              Port_n_name : mode data_type  
               );  
     END entity_name;  