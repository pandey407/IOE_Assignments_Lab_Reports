CONFIGURATION configuration_name OF entity_name IS  
FOR architecture_name  
  FOR instance_label : component_name  
     USE ENTITY library_name.entity_name(architecture_name);  
END FOR;  
END FOR;  
END [CONFIGURATION] [configuration_name];  