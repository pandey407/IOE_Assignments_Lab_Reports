ARCHITECTURE architecture_name OF entity_name IS  
BEGIN  
   (concurrent statements )  
END architecture_name;  